module register_input(alu_result_bus, eip, ebp, esp);
input [7:0]alu_result_bus;
output [7:0]eip;
output [7:0]ebp;
output [7:0]esp;


endmodule
